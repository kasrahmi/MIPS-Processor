library verilog;
use verilog.vl_types.all;
entity dCache_vlg_vec_tst is
end dCache_vlg_vec_tst;
