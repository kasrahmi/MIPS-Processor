library verilog;
use verilog.vl_types.all;
entity iCache_vlg_vec_tst is
end iCache_vlg_vec_tst;
