library verilog;
use verilog.vl_types.all;
entity triBufferbit8_vlg_vec_tst is
end triBufferbit8_vlg_vec_tst;
