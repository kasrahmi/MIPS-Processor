library verilog;
use verilog.vl_types.all;
entity pc2edges_vlg_vec_tst is
end pc2edges_vlg_vec_tst;
